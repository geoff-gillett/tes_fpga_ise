library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity file_io_TB is
end entity file_io_TB;

architecture RTL of file_io_TB is
	
begin

process 

end architecture RTL;
